module cau8(SW, KEY, LEDR);
	input [9:9]SW;
	input [0:0]KEY; // t = SW9, clk = KEY0
	output [0:0]LEDR;   // q = LEDR
	
	FF_T(SW[9], KEY[0], LEDR[0]);
endmodule

module FF_T(t, clk, q);
	input t, clk;
	output q;
	wire m1, m2, d;
	
	and(m1, ~t, q);
	and(m2, t, ~q);
	or(d, m1, m2);
	FF_D(d, clk, q);
endmodule

module FF_D(d, clk, q);
	input d, clk;
	output reg q;
	
	always @(posedge clk)
		q <= d;
endmodule

