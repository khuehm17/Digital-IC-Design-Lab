library verilog;
use verilog.vl_types.all;
entity cau1_vlg_tst is
end cau1_vlg_tst;
