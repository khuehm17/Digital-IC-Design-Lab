library verilog;
use verilog.vl_types.all;
entity cau2_vlg_vec_tst is
end cau2_vlg_vec_tst;
