library verilog;
use verilog.vl_types.all;
entity cau5_vlg_vec_tst is
end cau5_vlg_vec_tst;
